`timescale 1ns / 1ps

module weights_rom(
    clk, addr, rom_out
    );
    input wire clk;
    input wire [7:0] addr;
    output wire [7:0] rom_out;
    
    reg [7:0] rom_reg = 0;
    assign rom_out = rom_reg;
     
    always @(negedge clk) begin
        case (addr) 
            8'b00000000 : rom_reg <= 8'b00111110;
            8'b00000001 : rom_reg <= 8'b00110110;
            8'b00000010 : rom_reg <= 8'b11110110;
            8'b00000011 : rom_reg <= 8'b01000001;
            8'b00000100 : rom_reg <= 8'b11000010;
            8'b00000101 : rom_reg <= 8'b01001010;
            8'b00000110 : rom_reg <= 8'b00011111;
            8'b00000111 : rom_reg <= 8'b00001101;
            8'b00001000 : rom_reg <= 8'b11101001;
            8'b00001001 : rom_reg <= 8'b11011000;
            8'b00001010 : rom_reg <= 8'b00010000;
            8'b00001011 : rom_reg <= 8'b11100010;
            8'b00001100 : rom_reg <= 8'b00011100;
            8'b00001101 : rom_reg <= 8'b00101001;
            8'b00001110 : rom_reg <= 8'b11101011;
            8'b00001111 : rom_reg <= 8'b00011110;
            8'b00010000 : rom_reg <= 8'b00101011;
            8'b00010001 : rom_reg <= 8'b11110110;
            8'b00010010 : rom_reg <= 8'b11111110;
            8'b00010011 : rom_reg <= 8'b11011111;
            8'b00010100 : rom_reg <= 8'b10110011;
            8'b00010101 : rom_reg <= 8'b10000110;
            8'b00010110 : rom_reg <= 8'b00010111;
            8'b00010111 : rom_reg <= 8'b00001111;
            8'b00011000 : rom_reg <= 8'b00011011;
            8'b00011001 : rom_reg <= 8'b11111110;
            8'b00011010 : rom_reg <= 8'b11101010;
            8'b00011011 : rom_reg <= 8'b00000000;
            8'b00011100 : rom_reg <= 8'b00000000;
            8'b00011101 : rom_reg <= 8'b00001000;
            8'b00011110 : rom_reg <= 8'b11111001;
            8'b00011111 : rom_reg <= 8'b00001000;
            8'b00100000 : rom_reg <= 8'b11111111;
            8'b00100001 : rom_reg <= 8'b11111000;
            8'b00100010 : rom_reg <= 8'b00001101;
            8'b00100011 : rom_reg <= 8'b11111111;
            8'b00100100 : rom_reg <= 8'b11111101;
            8'b00100101 : rom_reg <= 8'b00101101;
            8'b00100110 : rom_reg <= 8'b00001100;
            8'b00100111 : rom_reg <= 8'b00100011;
            8'b00101000 : rom_reg <= 8'b00000000;
            8'b00101001 : rom_reg <= 8'b00000110;
            8'b00101010 : rom_reg <= 8'b00100100;
            8'b00101011 : rom_reg <= 8'b00111000;
            8'b00101100 : rom_reg <= 8'b00000011;
            8'b00101101 : rom_reg <= 8'b00011101;
            8'b00101110 : rom_reg <= 8'b00000010;
            8'b00101111 : rom_reg <= 8'b00111010;
            8'b00110000 : rom_reg <= 8'b00110010;
            8'b00110001 : rom_reg <= 8'b11111000;
            8'b00110010 : rom_reg <= 8'b00010110;
            8'b00110011 : rom_reg <= 8'b00001100;
            8'b00110100 : rom_reg <= 8'b00000110;
            8'b00110101 : rom_reg <= 8'b00000000;
            8'b00110110 : rom_reg <= 8'b00001111;
            8'b00110111 : rom_reg <= 8'b01000111;
            8'b00111000 : rom_reg <= 8'b01000010;
            8'b00111001 : rom_reg <= 8'b00001111;
            8'b00111010 : rom_reg <= 8'b00110010;
            8'b00111011 : rom_reg <= 8'b00010011;
            8'b00111100 : rom_reg <= 8'b00000111;
            8'b00111101 : rom_reg <= 8'b00011001;
            8'b00111110 : rom_reg <= 8'b11111110;
            8'b00111111 : rom_reg <= 8'b11100110;
            8'b01000000 : rom_reg <= 8'b11010001;
            8'b01000001 : rom_reg <= 8'b11100001;
            8'b01000010 : rom_reg <= 8'b11011011;
            8'b01000011 : rom_reg <= 8'b00000011;
            8'b01000100 : rom_reg <= 8'b11110011;
            8'b01000101 : rom_reg <= 8'b11001100;
            8'b01000110 : rom_reg <= 8'b11011011;
            8'b01000111 : rom_reg <= 8'b00100001;
            8'b01001000 : rom_reg <= 8'b00001110;
            8'b01001001 : rom_reg <= 8'b11111011;
            8'b01001010 : rom_reg <= 8'b00001011;
            8'b01001011 : rom_reg <= 8'b00000000;
            8'b01001100 : rom_reg <= 8'b00001101;
            8'b01001101 : rom_reg <= 8'b11101001;
            8'b01001110 : rom_reg <= 8'b11111111;
            8'b01001111 : rom_reg <= 8'b00010110;
            8'b01010000 : rom_reg <= 8'b00011011;
            8'b01010001 : rom_reg <= 8'b11110111;
            8'b01010010 : rom_reg <= 8'b11101010;
            8'b01010011 : rom_reg <= 8'b11101101;
            8'b01010100 : rom_reg <= 8'b11111000;
            8'b01010101 : rom_reg <= 8'b11101100;
            8'b01010110 : rom_reg <= 8'b00010000;
            8'b01010111 : rom_reg <= 8'b11010001;
            8'b01011000 : rom_reg <= 8'b00000001;
            8'b01011001 : rom_reg <= 8'b00000101;
            8'b01011010 : rom_reg <= 8'b11001111;


            default : rom_reg <= 8'b00000000;  
        endcase
    end
endmodule
