`timescale 1ns / 1ps
module tanh_lut #(parameter N=10, parameter Q=8) (
	input [N-1:0] addr,
	 input clk,
	 output signed [N-1:0] tanh_out
	);
reg signed [N-1:0] tanh_out_reg;
assign tanh_out = tanh_out_reg;

always @(negedge clk) begin
	case (addr)
		12'b0000000000 : tanh_out_reg <= 10'b0000000000;
		12'b0000000001 : tanh_out_reg <= 10'b0000000000;
		12'b0000000010 : tanh_out_reg <= 10'b0000000001;
		12'b0000000011 : tanh_out_reg <= 10'b0000000010;
		12'b0000000100 : tanh_out_reg <= 10'b0000000011;
		12'b0000000101 : tanh_out_reg <= 10'b0000000100;
		12'b0000000110 : tanh_out_reg <= 10'b0000000101;
		12'b0000000111 : tanh_out_reg <= 10'b0000000110;
		12'b0000001000 : tanh_out_reg <= 10'b0000000111;
		12'b0000001001 : tanh_out_reg <= 10'b0000001000;
		12'b0000001010 : tanh_out_reg <= 10'b0000001001;
		12'b0000001011 : tanh_out_reg <= 10'b0000001010;
		12'b0000001100 : tanh_out_reg <= 10'b0000001011;
		12'b0000001101 : tanh_out_reg <= 10'b0000001100;
		12'b0000001110 : tanh_out_reg <= 10'b0000001101;
		12'b0000001111 : tanh_out_reg <= 10'b0000001110;
		12'b0000010000 : tanh_out_reg <= 10'b0000001111;
		12'b0000010001 : tanh_out_reg <= 10'b0000010000;
		12'b0000010010 : tanh_out_reg <= 10'b0000010001;
		12'b0000010011 : tanh_out_reg <= 10'b0000010010;
		12'b0000010100 : tanh_out_reg <= 10'b0000010011;
		12'b0000010101 : tanh_out_reg <= 10'b0000010100;
		12'b0000010110 : tanh_out_reg <= 10'b0000010101;
		12'b0000010111 : tanh_out_reg <= 10'b0000010110;
		12'b0000011000 : tanh_out_reg <= 10'b0000010111;
		12'b0000011001 : tanh_out_reg <= 10'b0000011000;
		12'b0000011010 : tanh_out_reg <= 10'b0000011001;
		12'b0000011011 : tanh_out_reg <= 10'b0000011010;
		12'b0000011100 : tanh_out_reg <= 10'b0000011011;
		12'b0000011101 : tanh_out_reg <= 10'b0000011100;
		12'b0000011110 : tanh_out_reg <= 10'b0000011101;
		12'b0000011111 : tanh_out_reg <= 10'b0000011110;
		12'b0000100000 : tanh_out_reg <= 10'b0000011111;
		12'b0000100001 : tanh_out_reg <= 10'b0000100000;
		12'b0000100010 : tanh_out_reg <= 10'b0000100001;
		12'b0000100011 : tanh_out_reg <= 10'b0000100010;
		12'b0000100100 : tanh_out_reg <= 10'b0000100011;
		12'b0000100101 : tanh_out_reg <= 10'b0000100100;
		12'b0000100110 : tanh_out_reg <= 10'b0000100101;
		12'b0000100111 : tanh_out_reg <= 10'b0000100110;
		12'b0000101000 : tanh_out_reg <= 10'b0000100111;
		12'b0000101001 : tanh_out_reg <= 10'b0000101000;
		12'b0000101010 : tanh_out_reg <= 10'b0000101001;
		12'b0000101011 : tanh_out_reg <= 10'b0000101010;
		12'b0000101100 : tanh_out_reg <= 10'b0000101011;
		12'b0000101101 : tanh_out_reg <= 10'b0000101100;
		12'b0000101110 : tanh_out_reg <= 10'b0000101101;
		12'b0000101111 : tanh_out_reg <= 10'b0000101110;
		12'b0000110000 : tanh_out_reg <= 10'b0000101111;
		12'b0000110001 : tanh_out_reg <= 10'b0000110000;
		12'b0000110010 : tanh_out_reg <= 10'b0000110001;
		12'b0000110011 : tanh_out_reg <= 10'b0000110010;
		12'b0000110100 : tanh_out_reg <= 10'b0000110011;
		12'b0000110101 : tanh_out_reg <= 10'b0000110100;
		12'b0000110110 : tanh_out_reg <= 10'b0000110101;
		12'b0000110111 : tanh_out_reg <= 10'b0000110110;
		12'b0000111000 : tanh_out_reg <= 10'b0000110111;
		12'b0000111001 : tanh_out_reg <= 10'b0000111000;
		12'b0000111010 : tanh_out_reg <= 10'b0000111001;
		12'b0000111011 : tanh_out_reg <= 10'b0000111001;
		12'b0000111100 : tanh_out_reg <= 10'b0000111010;
		12'b0000111101 : tanh_out_reg <= 10'b0000111011;
		12'b0000111110 : tanh_out_reg <= 10'b0000111100;
		12'b0000111111 : tanh_out_reg <= 10'b0000111101;
		12'b0001000000 : tanh_out_reg <= 10'b0000111110;
		12'b0001000001 : tanh_out_reg <= 10'b0000111111;
		12'b0001000010 : tanh_out_reg <= 10'b0001000000;
		12'b0001000011 : tanh_out_reg <= 10'b0001000001;
		12'b0001000100 : tanh_out_reg <= 10'b0001000010;
		12'b0001000101 : tanh_out_reg <= 10'b0001000011;
		12'b0001000110 : tanh_out_reg <= 10'b0001000100;
		12'b0001000111 : tanh_out_reg <= 10'b0001000101;
		12'b0001001000 : tanh_out_reg <= 10'b0001000110;
		12'b0001001001 : tanh_out_reg <= 10'b0001000111;
		12'b0001001010 : tanh_out_reg <= 10'b0001001000;
		12'b0001001011 : tanh_out_reg <= 10'b0001001000;
		12'b0001001100 : tanh_out_reg <= 10'b0001001001;
		12'b0001001101 : tanh_out_reg <= 10'b0001001010;
		12'b0001001110 : tanh_out_reg <= 10'b0001001011;
		12'b0001001111 : tanh_out_reg <= 10'b0001001100;
		12'b0001010000 : tanh_out_reg <= 10'b0001001101;
		12'b0001010001 : tanh_out_reg <= 10'b0001001110;
		12'b0001010010 : tanh_out_reg <= 10'b0001001111;
		12'b0001010011 : tanh_out_reg <= 10'b0001010000;
		12'b0001010100 : tanh_out_reg <= 10'b0001010001;
		12'b0001010101 : tanh_out_reg <= 10'b0001010010;
		12'b0001010110 : tanh_out_reg <= 10'b0001010010;
		12'b0001010111 : tanh_out_reg <= 10'b0001010011;
		12'b0001011000 : tanh_out_reg <= 10'b0001010100;
		12'b0001011001 : tanh_out_reg <= 10'b0001010101;
		12'b0001011010 : tanh_out_reg <= 10'b0001010110;
		12'b0001011011 : tanh_out_reg <= 10'b0001010111;
		12'b0001011100 : tanh_out_reg <= 10'b0001011000;
		12'b0001011101 : tanh_out_reg <= 10'b0001011001;
		12'b0001011110 : tanh_out_reg <= 10'b0001011001;
		12'b0001011111 : tanh_out_reg <= 10'b0001011010;
		12'b0001100000 : tanh_out_reg <= 10'b0001011011;
		12'b0001100001 : tanh_out_reg <= 10'b0001011100;
		12'b0001100010 : tanh_out_reg <= 10'b0001011101;
		12'b0001100011 : tanh_out_reg <= 10'b0001011110;
		12'b0001100100 : tanh_out_reg <= 10'b0001011111;
		12'b0001100101 : tanh_out_reg <= 10'b0001100000;
		12'b0001100110 : tanh_out_reg <= 10'b0001100000;
		12'b0001100111 : tanh_out_reg <= 10'b0001100001;
		12'b0001101000 : tanh_out_reg <= 10'b0001100010;
		12'b0001101001 : tanh_out_reg <= 10'b0001100011;
		12'b0001101010 : tanh_out_reg <= 10'b0001100100;
		12'b0001101011 : tanh_out_reg <= 10'b0001100101;
		12'b0001101100 : tanh_out_reg <= 10'b0001100110;
		12'b0001101101 : tanh_out_reg <= 10'b0001100110;
		12'b0001101110 : tanh_out_reg <= 10'b0001100111;
		12'b0001101111 : tanh_out_reg <= 10'b0001101000;
		12'b0001110000 : tanh_out_reg <= 10'b0001101001;
		12'b0001110001 : tanh_out_reg <= 10'b0001101010;
		12'b0001110010 : tanh_out_reg <= 10'b0001101011;
		12'b0001110011 : tanh_out_reg <= 10'b0001101011;
		12'b0001110100 : tanh_out_reg <= 10'b0001101100;
		12'b0001110101 : tanh_out_reg <= 10'b0001101101;
		12'b0001110110 : tanh_out_reg <= 10'b0001101110;
		12'b0001110111 : tanh_out_reg <= 10'b0001101111;
		12'b0001111000 : tanh_out_reg <= 10'b0001101111;
		12'b0001111001 : tanh_out_reg <= 10'b0001110000;
		12'b0001111010 : tanh_out_reg <= 10'b0001110001;
		12'b0001111011 : tanh_out_reg <= 10'b0001110010;
		12'b0001111100 : tanh_out_reg <= 10'b0001110011;
		12'b0001111101 : tanh_out_reg <= 10'b0001110011;
		12'b0001111110 : tanh_out_reg <= 10'b0001110100;
		12'b0001111111 : tanh_out_reg <= 10'b0001110101;
		12'b0010000000 : tanh_out_reg <= 10'b0001110110;
		12'b0010000001 : tanh_out_reg <= 10'b0001110111;
		12'b0010000010 : tanh_out_reg <= 10'b0001110111;
		12'b0010000011 : tanh_out_reg <= 10'b0001111000;
		12'b0010000100 : tanh_out_reg <= 10'b0001111001;
		12'b0010000101 : tanh_out_reg <= 10'b0001111010;
		12'b0010000110 : tanh_out_reg <= 10'b0001111010;
		12'b0010000111 : tanh_out_reg <= 10'b0001111011;
		12'b0010001000 : tanh_out_reg <= 10'b0001111100;
		12'b0010001001 : tanh_out_reg <= 10'b0001111101;
		12'b0010001010 : tanh_out_reg <= 10'b0001111110;
		12'b0010001011 : tanh_out_reg <= 10'b0001111110;
		12'b0010001100 : tanh_out_reg <= 10'b0001111111;
		12'b0010001101 : tanh_out_reg <= 10'b0010000000;
		12'b0010001110 : tanh_out_reg <= 10'b0010000001;
		12'b0010001111 : tanh_out_reg <= 10'b0010000001;
		12'b0010010000 : tanh_out_reg <= 10'b0010000010;
		12'b0010010001 : tanh_out_reg <= 10'b0010000011;
		12'b0010010010 : tanh_out_reg <= 10'b0010000011;
		12'b0010010011 : tanh_out_reg <= 10'b0010000100;
		12'b0010010100 : tanh_out_reg <= 10'b0010000101;
		12'b0010010101 : tanh_out_reg <= 10'b0010000110;
		12'b0010010110 : tanh_out_reg <= 10'b0010000110;
		12'b0010010111 : tanh_out_reg <= 10'b0010000111;
		12'b0010011000 : tanh_out_reg <= 10'b0010001000;
		12'b0010011001 : tanh_out_reg <= 10'b0010001001;
		12'b0010011010 : tanh_out_reg <= 10'b0010001001;
		12'b0010011011 : tanh_out_reg <= 10'b0010001010;
		12'b0010011100 : tanh_out_reg <= 10'b0010001011;
		12'b0010011101 : tanh_out_reg <= 10'b0010001011;
		12'b0010011110 : tanh_out_reg <= 10'b0010001100;
		12'b0010011111 : tanh_out_reg <= 10'b0010001101;
		12'b0010100000 : tanh_out_reg <= 10'b0010001101;
		12'b0010100001 : tanh_out_reg <= 10'b0010001110;
		12'b0010100010 : tanh_out_reg <= 10'b0010001111;
		12'b0010100011 : tanh_out_reg <= 10'b0010010000;
		12'b0010100100 : tanh_out_reg <= 10'b0010010000;
		12'b0010100101 : tanh_out_reg <= 10'b0010010001;
		12'b0010100110 : tanh_out_reg <= 10'b0010010010;
		12'b0010100111 : tanh_out_reg <= 10'b0010010010;
		12'b0010101000 : tanh_out_reg <= 10'b0010010011;
		12'b0010101001 : tanh_out_reg <= 10'b0010010100;
		12'b0010101010 : tanh_out_reg <= 10'b0010010100;
		12'b0010101011 : tanh_out_reg <= 10'b0010010101;
		12'b0010101100 : tanh_out_reg <= 10'b0010010110;
		12'b0010101101 : tanh_out_reg <= 10'b0010010110;
		12'b0010101110 : tanh_out_reg <= 10'b0010010111;
		12'b0010101111 : tanh_out_reg <= 10'b0010011000;
		12'b0010110000 : tanh_out_reg <= 10'b0010011000;
		12'b0010110001 : tanh_out_reg <= 10'b0010011001;
		12'b0010110010 : tanh_out_reg <= 10'b0010011001;
		12'b0010110011 : tanh_out_reg <= 10'b0010011010;
		12'b0010110100 : tanh_out_reg <= 10'b0010011011;
		12'b0010110101 : tanh_out_reg <= 10'b0010011011;
		12'b0010110110 : tanh_out_reg <= 10'b0010011100;
		12'b0010110111 : tanh_out_reg <= 10'b0010011101;
		12'b0010111000 : tanh_out_reg <= 10'b0010011101;
		12'b0010111001 : tanh_out_reg <= 10'b0010011110;
		12'b0010111010 : tanh_out_reg <= 10'b0010011110;
		12'b0010111011 : tanh_out_reg <= 10'b0010011111;
		12'b0010111100 : tanh_out_reg <= 10'b0010100000;
		12'b0010111101 : tanh_out_reg <= 10'b0010100000;
		12'b0010111110 : tanh_out_reg <= 10'b0010100001;
		12'b0010111111 : tanh_out_reg <= 10'b0010100010;
		12'b0011000000 : tanh_out_reg <= 10'b0010100010;
		12'b0011000001 : tanh_out_reg <= 10'b0010100011;
		12'b0011000010 : tanh_out_reg <= 10'b0010100011;
		12'b0011000011 : tanh_out_reg <= 10'b0010100100;
		12'b0011000100 : tanh_out_reg <= 10'b0010100100;
		12'b0011000101 : tanh_out_reg <= 10'b0010100101;
		12'b0011000110 : tanh_out_reg <= 10'b0010100110;
		12'b0011000111 : tanh_out_reg <= 10'b0010100110;
		12'b0011001000 : tanh_out_reg <= 10'b0010100111;
		12'b0011001001 : tanh_out_reg <= 10'b0010100111;
		12'b0011001010 : tanh_out_reg <= 10'b0010101000;
		12'b0011001011 : tanh_out_reg <= 10'b0010101000;
		12'b0011001100 : tanh_out_reg <= 10'b0010101001;
		12'b0011001101 : tanh_out_reg <= 10'b0010101010;
		12'b0011001110 : tanh_out_reg <= 10'b0010101010;
		12'b0011001111 : tanh_out_reg <= 10'b0010101011;
		12'b0011010000 : tanh_out_reg <= 10'b0010101011;
		12'b0011010001 : tanh_out_reg <= 10'b0010101100;
		12'b0011010010 : tanh_out_reg <= 10'b0010101100;
		12'b0011010011 : tanh_out_reg <= 10'b0010101101;
		12'b0011010100 : tanh_out_reg <= 10'b0010101101;
		12'b0011010101 : tanh_out_reg <= 10'b0010101110;
		12'b0011010110 : tanh_out_reg <= 10'b0010101111;
		12'b0011010111 : tanh_out_reg <= 10'b0010101111;
		12'b0011011000 : tanh_out_reg <= 10'b0010110000;
		12'b0011011001 : tanh_out_reg <= 10'b0010110000;
		12'b0011011010 : tanh_out_reg <= 10'b0010110001;
		12'b0011011011 : tanh_out_reg <= 10'b0010110001;
		12'b0011011100 : tanh_out_reg <= 10'b0010110010;
		12'b0011011101 : tanh_out_reg <= 10'b0010110010;
		12'b0011011110 : tanh_out_reg <= 10'b0010110011;
		12'b0011011111 : tanh_out_reg <= 10'b0010110011;
		12'b0011100000 : tanh_out_reg <= 10'b0010110100;
		12'b0011100001 : tanh_out_reg <= 10'b0010110100;
		12'b0011100010 : tanh_out_reg <= 10'b0010110101;
		12'b0011100011 : tanh_out_reg <= 10'b0010110101;
		12'b0011100100 : tanh_out_reg <= 10'b0010110110;
		12'b0011100101 : tanh_out_reg <= 10'b0010110110;
		12'b0011100110 : tanh_out_reg <= 10'b0010110111;
		12'b0011100111 : tanh_out_reg <= 10'b0010110111;
		12'b0011101000 : tanh_out_reg <= 10'b0010111000;
		12'b0011101001 : tanh_out_reg <= 10'b0010111000;
		12'b0011101010 : tanh_out_reg <= 10'b0010111001;
		12'b0011101011 : tanh_out_reg <= 10'b0010111001;
		12'b0011101100 : tanh_out_reg <= 10'b0010111010;
		12'b0011101101 : tanh_out_reg <= 10'b0010111010;
		12'b0011101110 : tanh_out_reg <= 10'b0010111010;
		12'b0011101111 : tanh_out_reg <= 10'b0010111011;
		12'b0011110000 : tanh_out_reg <= 10'b0010111011;
		12'b0011110001 : tanh_out_reg <= 10'b0010111100;
		12'b0011110010 : tanh_out_reg <= 10'b0010111100;
		12'b0011110011 : tanh_out_reg <= 10'b0010111101;
		12'b0011110100 : tanh_out_reg <= 10'b0010111101;
		12'b0011110101 : tanh_out_reg <= 10'b0010111110;
		12'b0011110110 : tanh_out_reg <= 10'b0010111110;
		12'b0011110111 : tanh_out_reg <= 10'b0010111111;
		12'b0011111000 : tanh_out_reg <= 10'b0010111111;
		12'b0011111001 : tanh_out_reg <= 10'b0010111111;
		12'b0011111010 : tanh_out_reg <= 10'b0011000000;
		12'b0011111011 : tanh_out_reg <= 10'b0011000000;
		12'b0011111100 : tanh_out_reg <= 10'b0011000001;
		12'b0011111101 : tanh_out_reg <= 10'b0011000001;
		12'b0011111110 : tanh_out_reg <= 10'b0011000010;
		12'b0011111111 : tanh_out_reg <= 10'b0011000010;
		12'b0100000000 : tanh_out_reg <= 10'b0011000010;
		12'b0100000001 : tanh_out_reg <= 10'b0011000011;
		12'b0100000010 : tanh_out_reg <= 10'b0011000011;
		12'b0100000011 : tanh_out_reg <= 10'b0011000100;
		12'b0100000100 : tanh_out_reg <= 10'b0011000100;
		12'b0100000101 : tanh_out_reg <= 10'b0011000101;
		12'b0100000110 : tanh_out_reg <= 10'b0011000101;
		12'b0100000111 : tanh_out_reg <= 10'b0011000101;
		12'b0100001000 : tanh_out_reg <= 10'b0011000110;
		12'b0100001001 : tanh_out_reg <= 10'b0011000110;
		12'b0100001010 : tanh_out_reg <= 10'b0011000111;
		12'b0100001011 : tanh_out_reg <= 10'b0011000111;
		12'b0100001100 : tanh_out_reg <= 10'b0011000111;
		12'b0100001101 : tanh_out_reg <= 10'b0011001000;
		12'b0100001110 : tanh_out_reg <= 10'b0011001000;
		12'b0100001111 : tanh_out_reg <= 10'b0011001000;
		12'b0100010000 : tanh_out_reg <= 10'b0011001001;
		12'b0100010001 : tanh_out_reg <= 10'b0011001001;
		12'b0100010010 : tanh_out_reg <= 10'b0011001010;
		12'b0100010011 : tanh_out_reg <= 10'b0011001010;
		12'b0100010100 : tanh_out_reg <= 10'b0011001010;
		12'b0100010101 : tanh_out_reg <= 10'b0011001011;
		12'b0100010110 : tanh_out_reg <= 10'b0011001011;
		12'b0100010111 : tanh_out_reg <= 10'b0011001011;
		12'b0100011000 : tanh_out_reg <= 10'b0011001100;
		12'b0100011001 : tanh_out_reg <= 10'b0011001100;
		12'b0100011010 : tanh_out_reg <= 10'b0011001101;
		12'b0100011011 : tanh_out_reg <= 10'b0011001101;
		12'b0100011100 : tanh_out_reg <= 10'b0011001101;
		12'b0100011101 : tanh_out_reg <= 10'b0011001110;
		12'b0100011110 : tanh_out_reg <= 10'b0011001110;
		12'b0100011111 : tanh_out_reg <= 10'b0011001110;
		12'b0100100000 : tanh_out_reg <= 10'b0011001111;
		12'b0100100001 : tanh_out_reg <= 10'b0011001111;
		12'b0100100010 : tanh_out_reg <= 10'b0011001111;
		12'b0100100011 : tanh_out_reg <= 10'b0011010000;
		12'b0100100100 : tanh_out_reg <= 10'b0011010000;
		12'b0100100101 : tanh_out_reg <= 10'b0011010000;
		12'b0100100110 : tanh_out_reg <= 10'b0011010001;
		12'b0100100111 : tanh_out_reg <= 10'b0011010001;
		12'b0100101000 : tanh_out_reg <= 10'b0011010001;
		12'b0100101001 : tanh_out_reg <= 10'b0011010010;
		12'b0100101010 : tanh_out_reg <= 10'b0011010010;
		12'b0100101011 : tanh_out_reg <= 10'b0011010010;
		12'b0100101100 : tanh_out_reg <= 10'b0011010011;
		12'b0100101101 : tanh_out_reg <= 10'b0011010011;
		12'b0100101110 : tanh_out_reg <= 10'b0011010011;
		12'b0100101111 : tanh_out_reg <= 10'b0011010100;
		12'b0100110000 : tanh_out_reg <= 10'b0011010100;
		12'b0100110001 : tanh_out_reg <= 10'b0011010100;
		12'b0100110010 : tanh_out_reg <= 10'b0011010101;
		12'b0100110011 : tanh_out_reg <= 10'b0011010101;
		12'b0100110100 : tanh_out_reg <= 10'b0011010101;
		12'b0100110101 : tanh_out_reg <= 10'b0011010101;
		12'b0100110110 : tanh_out_reg <= 10'b0011010110;
		12'b0100110111 : tanh_out_reg <= 10'b0011010110;
		12'b0100111000 : tanh_out_reg <= 10'b0011010110;
		12'b0100111001 : tanh_out_reg <= 10'b0011010111;
		12'b0100111010 : tanh_out_reg <= 10'b0011010111;
		12'b0100111011 : tanh_out_reg <= 10'b0011010111;
		12'b0100111100 : tanh_out_reg <= 10'b0011011000;
		12'b0100111101 : tanh_out_reg <= 10'b0011011000;
		12'b0100111110 : tanh_out_reg <= 10'b0011011000;
		12'b0100111111 : tanh_out_reg <= 10'b0011011000;
		12'b0101000000 : tanh_out_reg <= 10'b0011011001;
		12'b0101000001 : tanh_out_reg <= 10'b0011011001;
		12'b0101000010 : tanh_out_reg <= 10'b0011011001;
		12'b0101000011 : tanh_out_reg <= 10'b0011011001;
		12'b0101000100 : tanh_out_reg <= 10'b0011011010;
		12'b0101000101 : tanh_out_reg <= 10'b0011011010;
		12'b0101000110 : tanh_out_reg <= 10'b0011011010;
		12'b0101000111 : tanh_out_reg <= 10'b0011011011;
		12'b0101001000 : tanh_out_reg <= 10'b0011011011;
		12'b0101001001 : tanh_out_reg <= 10'b0011011011;
		12'b0101001010 : tanh_out_reg <= 10'b0011011011;
		12'b0101001011 : tanh_out_reg <= 10'b0011011100;
		12'b0101001100 : tanh_out_reg <= 10'b0011011100;
		12'b0101001101 : tanh_out_reg <= 10'b0011011100;
		12'b0101001110 : tanh_out_reg <= 10'b0011011100;
		12'b0101001111 : tanh_out_reg <= 10'b0011011101;
		12'b0101010000 : tanh_out_reg <= 10'b0011011101;
		12'b0101010001 : tanh_out_reg <= 10'b0011011101;
		12'b0101010010 : tanh_out_reg <= 10'b0011011101;
		12'b0101010011 : tanh_out_reg <= 10'b0011011110;
		12'b0101010100 : tanh_out_reg <= 10'b0011011110;
		12'b0101010101 : tanh_out_reg <= 10'b0011011110;
		12'b0101010110 : tanh_out_reg <= 10'b0011011110;
		12'b0101010111 : tanh_out_reg <= 10'b0011011111;
		12'b0101011000 : tanh_out_reg <= 10'b0011011111;
		12'b0101011001 : tanh_out_reg <= 10'b0011011111;
		12'b0101011010 : tanh_out_reg <= 10'b0011011111;
		12'b0101011011 : tanh_out_reg <= 10'b0011100000;
		12'b0101011100 : tanh_out_reg <= 10'b0011100000;
		12'b0101011101 : tanh_out_reg <= 10'b0011100000;
		12'b0101011110 : tanh_out_reg <= 10'b0011100000;
		12'b0101011111 : tanh_out_reg <= 10'b0011100001;
		12'b0101100000 : tanh_out_reg <= 10'b0011100001;
		12'b0101100001 : tanh_out_reg <= 10'b0011100001;
		12'b0101100010 : tanh_out_reg <= 10'b0011100001;
		12'b0101100011 : tanh_out_reg <= 10'b0011100001;
		12'b0101100100 : tanh_out_reg <= 10'b0011100010;
		12'b0101100101 : tanh_out_reg <= 10'b0011100010;
		12'b0101100110 : tanh_out_reg <= 10'b0011100010;
		12'b0101100111 : tanh_out_reg <= 10'b0011100010;
		12'b0101101000 : tanh_out_reg <= 10'b0011100010;
		12'b0101101001 : tanh_out_reg <= 10'b0011100011;
		12'b0101101010 : tanh_out_reg <= 10'b0011100011;
		12'b0101101011 : tanh_out_reg <= 10'b0011100011;
		12'b0101101100 : tanh_out_reg <= 10'b0011100011;
		12'b0101101101 : tanh_out_reg <= 10'b0011100100;
		12'b0101101110 : tanh_out_reg <= 10'b0011100100;
		12'b0101101111 : tanh_out_reg <= 10'b0011100100;
		12'b0101110000 : tanh_out_reg <= 10'b0011100100;
		12'b0101110001 : tanh_out_reg <= 10'b0011100100;
		12'b0101110010 : tanh_out_reg <= 10'b0011100101;
		12'b0101110011 : tanh_out_reg <= 10'b0011100101;
		12'b0101110100 : tanh_out_reg <= 10'b0011100101;
		12'b0101110101 : tanh_out_reg <= 10'b0011100101;
		12'b0101110110 : tanh_out_reg <= 10'b0011100101;
		12'b0101110111 : tanh_out_reg <= 10'b0011100110;
		12'b0101111000 : tanh_out_reg <= 10'b0011100110;
		12'b0101111001 : tanh_out_reg <= 10'b0011100110;
		12'b0101111010 : tanh_out_reg <= 10'b0011100110;
		12'b0101111011 : tanh_out_reg <= 10'b0011100110;
		12'b0101111100 : tanh_out_reg <= 10'b0011100110;
		12'b0101111101 : tanh_out_reg <= 10'b0011100111;
		12'b0101111110 : tanh_out_reg <= 10'b0011100111;
		12'b0101111111 : tanh_out_reg <= 10'b0011100111;
		12'b0110000000 : tanh_out_reg <= 10'b0011100111;
		12'b0110000001 : tanh_out_reg <= 10'b0011100111;
		12'b0110000010 : tanh_out_reg <= 10'b0011101000;
		12'b0110000011 : tanh_out_reg <= 10'b0011101000;
		12'b0110000100 : tanh_out_reg <= 10'b0011101000;
		12'b0110000101 : tanh_out_reg <= 10'b0011101000;
		12'b0110000110 : tanh_out_reg <= 10'b0011101000;
		12'b0110000111 : tanh_out_reg <= 10'b0011101000;
		12'b0110001000 : tanh_out_reg <= 10'b0011101001;
		12'b0110001001 : tanh_out_reg <= 10'b0011101001;
		12'b0110001010 : tanh_out_reg <= 10'b0011101001;
		12'b0110001011 : tanh_out_reg <= 10'b0011101001;
		12'b0110001100 : tanh_out_reg <= 10'b0011101001;
		12'b0110001101 : tanh_out_reg <= 10'b0011101001;
		12'b0110001110 : tanh_out_reg <= 10'b0011101010;
		12'b0110001111 : tanh_out_reg <= 10'b0011101010;
		12'b0110010000 : tanh_out_reg <= 10'b0011101010;
		12'b0110010001 : tanh_out_reg <= 10'b0011101010;
		12'b0110010010 : tanh_out_reg <= 10'b0011101010;
		12'b0110010011 : tanh_out_reg <= 10'b0011101010;
		12'b0110010100 : tanh_out_reg <= 10'b0011101011;
		12'b0110010101 : tanh_out_reg <= 10'b0011101011;
		12'b0110010110 : tanh_out_reg <= 10'b0011101011;
		12'b0110010111 : tanh_out_reg <= 10'b0011101011;
		12'b0110011000 : tanh_out_reg <= 10'b0011101011;
		12'b0110011001 : tanh_out_reg <= 10'b0011101011;
		12'b0110011010 : tanh_out_reg <= 10'b0011101100;
		12'b0110011011 : tanh_out_reg <= 10'b0011101100;
		12'b0110011100 : tanh_out_reg <= 10'b0011101100;
		12'b0110011101 : tanh_out_reg <= 10'b0011101100;
		12'b0110011110 : tanh_out_reg <= 10'b0011101100;
		12'b0110011111 : tanh_out_reg <= 10'b0011101100;
		12'b0110100000 : tanh_out_reg <= 10'b0011101100;
		12'b0110100001 : tanh_out_reg <= 10'b0011101101;
		12'b0110100010 : tanh_out_reg <= 10'b0011101101;
		12'b0110100011 : tanh_out_reg <= 10'b0011101101;
		12'b0110100100 : tanh_out_reg <= 10'b0011101101;
		12'b0110100101 : tanh_out_reg <= 10'b0011101101;
		12'b0110100110 : tanh_out_reg <= 10'b0011101101;
		12'b0110100111 : tanh_out_reg <= 10'b0011101101;
		12'b0110101000 : tanh_out_reg <= 10'b0011101110;
		12'b0110101001 : tanh_out_reg <= 10'b0011101110;
		12'b0110101010 : tanh_out_reg <= 10'b0011101110;
		12'b0110101011 : tanh_out_reg <= 10'b0011101110;
		12'b0110101100 : tanh_out_reg <= 10'b0011101110;
		12'b0110101101 : tanh_out_reg <= 10'b0011101110;
		12'b0110101110 : tanh_out_reg <= 10'b0011101110;
		12'b0110101111 : tanh_out_reg <= 10'b0011101110;
		12'b0110110000 : tanh_out_reg <= 10'b0011101111;
		12'b0110110001 : tanh_out_reg <= 10'b0011101111;
		12'b0110110010 : tanh_out_reg <= 10'b0011101111;
		12'b0110110011 : tanh_out_reg <= 10'b0011101111;
		12'b0110110100 : tanh_out_reg <= 10'b0011101111;
		12'b0110110101 : tanh_out_reg <= 10'b0011101111;
		12'b0110110110 : tanh_out_reg <= 10'b0011101111;
		12'b0110110111 : tanh_out_reg <= 10'b0011101111;
		12'b0110111000 : tanh_out_reg <= 10'b0011110000;
		12'b0110111001 : tanh_out_reg <= 10'b0011110000;
		12'b0110111010 : tanh_out_reg <= 10'b0011110000;
		12'b0110111011 : tanh_out_reg <= 10'b0011110000;
		12'b0110111100 : tanh_out_reg <= 10'b0011110000;
		12'b0110111101 : tanh_out_reg <= 10'b0011110000;
		12'b0110111110 : tanh_out_reg <= 10'b0011110000;
		12'b0110111111 : tanh_out_reg <= 10'b0011110000;
		12'b0111000000 : tanh_out_reg <= 10'b0011110000;
		12'b0111000001 : tanh_out_reg <= 10'b0011110001;
		12'b0111000010 : tanh_out_reg <= 10'b0011110001;
		12'b0111000011 : tanh_out_reg <= 10'b0011110001;
		12'b0111000100 : tanh_out_reg <= 10'b0011110001;
		12'b0111000101 : tanh_out_reg <= 10'b0011110001;
		12'b0111000110 : tanh_out_reg <= 10'b0011110001;
		12'b0111000111 : tanh_out_reg <= 10'b0011110001;
		12'b0111001000 : tanh_out_reg <= 10'b0011110001;
		12'b0111001001 : tanh_out_reg <= 10'b0011110001;
		12'b0111001010 : tanh_out_reg <= 10'b0011110010;
		12'b0111001011 : tanh_out_reg <= 10'b0011110010;
		12'b0111001100 : tanh_out_reg <= 10'b0011110010;
		12'b0111001101 : tanh_out_reg <= 10'b0011110010;
		12'b0111001110 : tanh_out_reg <= 10'b0011110010;
		12'b0111001111 : tanh_out_reg <= 10'b0011110010;
		12'b0111010000 : tanh_out_reg <= 10'b0011110010;
		12'b0111010001 : tanh_out_reg <= 10'b0011110010;
		12'b0111010010 : tanh_out_reg <= 10'b0011110010;
		12'b0111010011 : tanh_out_reg <= 10'b0011110011;
		12'b0111010100 : tanh_out_reg <= 10'b0011110011;
		12'b0111010101 : tanh_out_reg <= 10'b0011110011;
		12'b0111010110 : tanh_out_reg <= 10'b0011110011;
		12'b0111010111 : tanh_out_reg <= 10'b0011110011;
		12'b0111011000 : tanh_out_reg <= 10'b0011110011;
		12'b0111011001 : tanh_out_reg <= 10'b0011110011;
		12'b0111011010 : tanh_out_reg <= 10'b0011110011;
		12'b0111011011 : tanh_out_reg <= 10'b0011110011;
		12'b0111011100 : tanh_out_reg <= 10'b0011110011;
		12'b0111011101 : tanh_out_reg <= 10'b0011110011;
		12'b0111011110 : tanh_out_reg <= 10'b0011110100;
		12'b0111011111 : tanh_out_reg <= 10'b0011110100;
		12'b0111100000 : tanh_out_reg <= 10'b0011110100;
		12'b0111100001 : tanh_out_reg <= 10'b0011110100;
		12'b0111100010 : tanh_out_reg <= 10'b0011110100;
		12'b0111100011 : tanh_out_reg <= 10'b0011110100;
		12'b0111100100 : tanh_out_reg <= 10'b0011110100;
		12'b0111100101 : tanh_out_reg <= 10'b0011110100;
		12'b0111100110 : tanh_out_reg <= 10'b0011110100;
		12'b0111100111 : tanh_out_reg <= 10'b0011110100;
		12'b0111101000 : tanh_out_reg <= 10'b0011110100;
		12'b0111101001 : tanh_out_reg <= 10'b0011110101;
		12'b0111101010 : tanh_out_reg <= 10'b0011110101;
		12'b0111101011 : tanh_out_reg <= 10'b0011110101;
		12'b0111101100 : tanh_out_reg <= 10'b0011110101;
		12'b0111101101 : tanh_out_reg <= 10'b0011110101;
		12'b0111101110 : tanh_out_reg <= 10'b0011110101;
		12'b0111101111 : tanh_out_reg <= 10'b0011110101;
		12'b0111110000 : tanh_out_reg <= 10'b0011110101;
		12'b0111110001 : tanh_out_reg <= 10'b0011110101;
		12'b0111110010 : tanh_out_reg <= 10'b0011110101;
		12'b0111110011 : tanh_out_reg <= 10'b0011110101;
		12'b0111110100 : tanh_out_reg <= 10'b0011110101;
		12'b0111110101 : tanh_out_reg <= 10'b0011110101;
		12'b0111110110 : tanh_out_reg <= 10'b0011110110;
		12'b0111110111 : tanh_out_reg <= 10'b0011110110;
		12'b0111111000 : tanh_out_reg <= 10'b0011110110;
		12'b0111111001 : tanh_out_reg <= 10'b0011110110;
		12'b0111111010 : tanh_out_reg <= 10'b0011110110;
		12'b0111111011 : tanh_out_reg <= 10'b0011110110;
		12'b0111111100 : tanh_out_reg <= 10'b0011110110;
		12'b0111111101 : tanh_out_reg <= 10'b0011110110;
		12'b0111111110 : tanh_out_reg <= 10'b0011110110;
		12'b0111111111 : tanh_out_reg <= 10'b0011110110;
		12'b1000000000 : tanh_out_reg <= 10'b1100001010;
		12'b1000000001 : tanh_out_reg <= 10'b1100001010;
		12'b1000000010 : tanh_out_reg <= 10'b1100001010;
		12'b1000000011 : tanh_out_reg <= 10'b1100001010;
		12'b1000000100 : tanh_out_reg <= 10'b1100001010;
		12'b1000000101 : tanh_out_reg <= 10'b1100001010;
		12'b1000000110 : tanh_out_reg <= 10'b1100001010;
		12'b1000000111 : tanh_out_reg <= 10'b1100001010;
		12'b1000001000 : tanh_out_reg <= 10'b1100001010;
		12'b1000001001 : tanh_out_reg <= 10'b1100001010;
		12'b1000001010 : tanh_out_reg <= 10'b1100001010;
		12'b1000001011 : tanh_out_reg <= 10'b1100001011;
		12'b1000001100 : tanh_out_reg <= 10'b1100001011;
		12'b1000001101 : tanh_out_reg <= 10'b1100001011;
		12'b1000001110 : tanh_out_reg <= 10'b1100001011;
		12'b1000001111 : tanh_out_reg <= 10'b1100001011;
		12'b1000010000 : tanh_out_reg <= 10'b1100001011;
		12'b1000010001 : tanh_out_reg <= 10'b1100001011;
		12'b1000010010 : tanh_out_reg <= 10'b1100001011;
		12'b1000010011 : tanh_out_reg <= 10'b1100001011;
		12'b1000010100 : tanh_out_reg <= 10'b1100001011;
		12'b1000010101 : tanh_out_reg <= 10'b1100001011;
		12'b1000010110 : tanh_out_reg <= 10'b1100001011;
		12'b1000010111 : tanh_out_reg <= 10'b1100001011;
		12'b1000011000 : tanh_out_reg <= 10'b1100001100;
		12'b1000011001 : tanh_out_reg <= 10'b1100001100;
		12'b1000011010 : tanh_out_reg <= 10'b1100001100;
		12'b1000011011 : tanh_out_reg <= 10'b1100001100;
		12'b1000011100 : tanh_out_reg <= 10'b1100001100;
		12'b1000011101 : tanh_out_reg <= 10'b1100001100;
		12'b1000011110 : tanh_out_reg <= 10'b1100001100;
		12'b1000011111 : tanh_out_reg <= 10'b1100001100;
		12'b1000100000 : tanh_out_reg <= 10'b1100001100;
		12'b1000100001 : tanh_out_reg <= 10'b1100001100;
		12'b1000100010 : tanh_out_reg <= 10'b1100001100;
		12'b1000100011 : tanh_out_reg <= 10'b1100001101;
		12'b1000100100 : tanh_out_reg <= 10'b1100001101;
		12'b1000100101 : tanh_out_reg <= 10'b1100001101;
		12'b1000100110 : tanh_out_reg <= 10'b1100001101;
		12'b1000100111 : tanh_out_reg <= 10'b1100001101;
		12'b1000101000 : tanh_out_reg <= 10'b1100001101;
		12'b1000101001 : tanh_out_reg <= 10'b1100001101;
		12'b1000101010 : tanh_out_reg <= 10'b1100001101;
		12'b1000101011 : tanh_out_reg <= 10'b1100001101;
		12'b1000101100 : tanh_out_reg <= 10'b1100001101;
		12'b1000101101 : tanh_out_reg <= 10'b1100001101;
		12'b1000101110 : tanh_out_reg <= 10'b1100001110;
		12'b1000101111 : tanh_out_reg <= 10'b1100001110;
		12'b1000110000 : tanh_out_reg <= 10'b1100001110;
		12'b1000110001 : tanh_out_reg <= 10'b1100001110;
		12'b1000110010 : tanh_out_reg <= 10'b1100001110;
		12'b1000110011 : tanh_out_reg <= 10'b1100001110;
		12'b1000110100 : tanh_out_reg <= 10'b1100001110;
		12'b1000110101 : tanh_out_reg <= 10'b1100001110;
		12'b1000110110 : tanh_out_reg <= 10'b1100001110;
		12'b1000110111 : tanh_out_reg <= 10'b1100001111;
		12'b1000111000 : tanh_out_reg <= 10'b1100001111;
		12'b1000111001 : tanh_out_reg <= 10'b1100001111;
		12'b1000111010 : tanh_out_reg <= 10'b1100001111;
		12'b1000111011 : tanh_out_reg <= 10'b1100001111;
		12'b1000111100 : tanh_out_reg <= 10'b1100001111;
		12'b1000111101 : tanh_out_reg <= 10'b1100001111;
		12'b1000111110 : tanh_out_reg <= 10'b1100001111;
		12'b1000111111 : tanh_out_reg <= 10'b1100001111;
		12'b1001000000 : tanh_out_reg <= 10'b1100010000;
		12'b1001000001 : tanh_out_reg <= 10'b1100010000;
		12'b1001000010 : tanh_out_reg <= 10'b1100010000;
		12'b1001000011 : tanh_out_reg <= 10'b1100010000;
		12'b1001000100 : tanh_out_reg <= 10'b1100010000;
		12'b1001000101 : tanh_out_reg <= 10'b1100010000;
		12'b1001000110 : tanh_out_reg <= 10'b1100010000;
		12'b1001000111 : tanh_out_reg <= 10'b1100010000;
		12'b1001001000 : tanh_out_reg <= 10'b1100010000;
		12'b1001001001 : tanh_out_reg <= 10'b1100010001;
		12'b1001001010 : tanh_out_reg <= 10'b1100010001;
		12'b1001001011 : tanh_out_reg <= 10'b1100010001;
		12'b1001001100 : tanh_out_reg <= 10'b1100010001;
		12'b1001001101 : tanh_out_reg <= 10'b1100010001;
		12'b1001001110 : tanh_out_reg <= 10'b1100010001;
		12'b1001001111 : tanh_out_reg <= 10'b1100010001;
		12'b1001010000 : tanh_out_reg <= 10'b1100010001;
		12'b1001010001 : tanh_out_reg <= 10'b1100010010;
		12'b1001010010 : tanh_out_reg <= 10'b1100010010;
		12'b1001010011 : tanh_out_reg <= 10'b1100010010;
		12'b1001010100 : tanh_out_reg <= 10'b1100010010;
		12'b1001010101 : tanh_out_reg <= 10'b1100010010;
		12'b1001010110 : tanh_out_reg <= 10'b1100010010;
		12'b1001010111 : tanh_out_reg <= 10'b1100010010;
		12'b1001011000 : tanh_out_reg <= 10'b1100010010;
		12'b1001011001 : tanh_out_reg <= 10'b1100010011;
		12'b1001011010 : tanh_out_reg <= 10'b1100010011;
		12'b1001011011 : tanh_out_reg <= 10'b1100010011;
		12'b1001011100 : tanh_out_reg <= 10'b1100010011;
		12'b1001011101 : tanh_out_reg <= 10'b1100010011;
		12'b1001011110 : tanh_out_reg <= 10'b1100010011;
		12'b1001011111 : tanh_out_reg <= 10'b1100010011;
		12'b1001100000 : tanh_out_reg <= 10'b1100010100;
		12'b1001100001 : tanh_out_reg <= 10'b1100010100;
		12'b1001100010 : tanh_out_reg <= 10'b1100010100;
		12'b1001100011 : tanh_out_reg <= 10'b1100010100;
		12'b1001100100 : tanh_out_reg <= 10'b1100010100;
		12'b1001100101 : tanh_out_reg <= 10'b1100010100;
		12'b1001100110 : tanh_out_reg <= 10'b1100010100;
		12'b1001100111 : tanh_out_reg <= 10'b1100010101;
		12'b1001101000 : tanh_out_reg <= 10'b1100010101;
		12'b1001101001 : tanh_out_reg <= 10'b1100010101;
		12'b1001101010 : tanh_out_reg <= 10'b1100010101;
		12'b1001101011 : tanh_out_reg <= 10'b1100010101;
		12'b1001101100 : tanh_out_reg <= 10'b1100010101;
		12'b1001101101 : tanh_out_reg <= 10'b1100010110;
		12'b1001101110 : tanh_out_reg <= 10'b1100010110;
		12'b1001101111 : tanh_out_reg <= 10'b1100010110;
		12'b1001110000 : tanh_out_reg <= 10'b1100010110;
		12'b1001110001 : tanh_out_reg <= 10'b1100010110;
		12'b1001110010 : tanh_out_reg <= 10'b1100010110;
		12'b1001110011 : tanh_out_reg <= 10'b1100010111;
		12'b1001110100 : tanh_out_reg <= 10'b1100010111;
		12'b1001110101 : tanh_out_reg <= 10'b1100010111;
		12'b1001110110 : tanh_out_reg <= 10'b1100010111;
		12'b1001110111 : tanh_out_reg <= 10'b1100010111;
		12'b1001111000 : tanh_out_reg <= 10'b1100010111;
		12'b1001111001 : tanh_out_reg <= 10'b1100011000;
		12'b1001111010 : tanh_out_reg <= 10'b1100011000;
		12'b1001111011 : tanh_out_reg <= 10'b1100011000;
		12'b1001111100 : tanh_out_reg <= 10'b1100011000;
		12'b1001111101 : tanh_out_reg <= 10'b1100011000;
		12'b1001111110 : tanh_out_reg <= 10'b1100011000;
		12'b1001111111 : tanh_out_reg <= 10'b1100011001;
		12'b1010000000 : tanh_out_reg <= 10'b1100011001;
		12'b1010000001 : tanh_out_reg <= 10'b1100011001;
		12'b1010000010 : tanh_out_reg <= 10'b1100011001;
		12'b1010000011 : tanh_out_reg <= 10'b1100011001;
		12'b1010000100 : tanh_out_reg <= 10'b1100011010;
		12'b1010000101 : tanh_out_reg <= 10'b1100011010;
		12'b1010000110 : tanh_out_reg <= 10'b1100011010;
		12'b1010000111 : tanh_out_reg <= 10'b1100011010;
		12'b1010001000 : tanh_out_reg <= 10'b1100011010;
		12'b1010001001 : tanh_out_reg <= 10'b1100011010;
		12'b1010001010 : tanh_out_reg <= 10'b1100011011;
		12'b1010001011 : tanh_out_reg <= 10'b1100011011;
		12'b1010001100 : tanh_out_reg <= 10'b1100011011;
		12'b1010001101 : tanh_out_reg <= 10'b1100011011;
		12'b1010001110 : tanh_out_reg <= 10'b1100011011;
		12'b1010001111 : tanh_out_reg <= 10'b1100011100;
		12'b1010010000 : tanh_out_reg <= 10'b1100011100;
		12'b1010010001 : tanh_out_reg <= 10'b1100011100;
		12'b1010010010 : tanh_out_reg <= 10'b1100011100;
		12'b1010010011 : tanh_out_reg <= 10'b1100011100;
		12'b1010010100 : tanh_out_reg <= 10'b1100011101;
		12'b1010010101 : tanh_out_reg <= 10'b1100011101;
		12'b1010010110 : tanh_out_reg <= 10'b1100011101;
		12'b1010010111 : tanh_out_reg <= 10'b1100011101;
		12'b1010011000 : tanh_out_reg <= 10'b1100011110;
		12'b1010011001 : tanh_out_reg <= 10'b1100011110;
		12'b1010011010 : tanh_out_reg <= 10'b1100011110;
		12'b1010011011 : tanh_out_reg <= 10'b1100011110;
		12'b1010011100 : tanh_out_reg <= 10'b1100011110;
		12'b1010011101 : tanh_out_reg <= 10'b1100011111;
		12'b1010011110 : tanh_out_reg <= 10'b1100011111;
		12'b1010011111 : tanh_out_reg <= 10'b1100011111;
		12'b1010100000 : tanh_out_reg <= 10'b1100011111;
		12'b1010100001 : tanh_out_reg <= 10'b1100011111;
		12'b1010100010 : tanh_out_reg <= 10'b1100100000;
		12'b1010100011 : tanh_out_reg <= 10'b1100100000;
		12'b1010100100 : tanh_out_reg <= 10'b1100100000;
		12'b1010100101 : tanh_out_reg <= 10'b1100100000;
		12'b1010100110 : tanh_out_reg <= 10'b1100100001;
		12'b1010100111 : tanh_out_reg <= 10'b1100100001;
		12'b1010101000 : tanh_out_reg <= 10'b1100100001;
		12'b1010101001 : tanh_out_reg <= 10'b1100100001;
		12'b1010101010 : tanh_out_reg <= 10'b1100100010;
		12'b1010101011 : tanh_out_reg <= 10'b1100100010;
		12'b1010101100 : tanh_out_reg <= 10'b1100100010;
		12'b1010101101 : tanh_out_reg <= 10'b1100100010;
		12'b1010101110 : tanh_out_reg <= 10'b1100100011;
		12'b1010101111 : tanh_out_reg <= 10'b1100100011;
		12'b1010110000 : tanh_out_reg <= 10'b1100100011;
		12'b1010110001 : tanh_out_reg <= 10'b1100100011;
		12'b1010110010 : tanh_out_reg <= 10'b1100100100;
		12'b1010110011 : tanh_out_reg <= 10'b1100100100;
		12'b1010110100 : tanh_out_reg <= 10'b1100100100;
		12'b1010110101 : tanh_out_reg <= 10'b1100100100;
		12'b1010110110 : tanh_out_reg <= 10'b1100100101;
		12'b1010110111 : tanh_out_reg <= 10'b1100100101;
		12'b1010111000 : tanh_out_reg <= 10'b1100100101;
		12'b1010111001 : tanh_out_reg <= 10'b1100100101;
		12'b1010111010 : tanh_out_reg <= 10'b1100100110;
		12'b1010111011 : tanh_out_reg <= 10'b1100100110;
		12'b1010111100 : tanh_out_reg <= 10'b1100100110;
		12'b1010111101 : tanh_out_reg <= 10'b1100100111;
		12'b1010111110 : tanh_out_reg <= 10'b1100100111;
		12'b1010111111 : tanh_out_reg <= 10'b1100100111;
		12'b1011000000 : tanh_out_reg <= 10'b1100100111;
		12'b1011000001 : tanh_out_reg <= 10'b1100101000;
		12'b1011000010 : tanh_out_reg <= 10'b1100101000;
		12'b1011000011 : tanh_out_reg <= 10'b1100101000;
		12'b1011000100 : tanh_out_reg <= 10'b1100101000;
		12'b1011000101 : tanh_out_reg <= 10'b1100101001;
		12'b1011000110 : tanh_out_reg <= 10'b1100101001;
		12'b1011000111 : tanh_out_reg <= 10'b1100101001;
		12'b1011001000 : tanh_out_reg <= 10'b1100101010;
		12'b1011001001 : tanh_out_reg <= 10'b1100101010;
		12'b1011001010 : tanh_out_reg <= 10'b1100101010;
		12'b1011001011 : tanh_out_reg <= 10'b1100101011;
		12'b1011001100 : tanh_out_reg <= 10'b1100101011;
		12'b1011001101 : tanh_out_reg <= 10'b1100101011;
		12'b1011001110 : tanh_out_reg <= 10'b1100101011;
		12'b1011001111 : tanh_out_reg <= 10'b1100101100;
		12'b1011010000 : tanh_out_reg <= 10'b1100101100;
		12'b1011010001 : tanh_out_reg <= 10'b1100101100;
		12'b1011010010 : tanh_out_reg <= 10'b1100101101;
		12'b1011010011 : tanh_out_reg <= 10'b1100101101;
		12'b1011010100 : tanh_out_reg <= 10'b1100101101;
		12'b1011010101 : tanh_out_reg <= 10'b1100101110;
		12'b1011010110 : tanh_out_reg <= 10'b1100101110;
		12'b1011010111 : tanh_out_reg <= 10'b1100101110;
		12'b1011011000 : tanh_out_reg <= 10'b1100101111;
		12'b1011011001 : tanh_out_reg <= 10'b1100101111;
		12'b1011011010 : tanh_out_reg <= 10'b1100101111;
		12'b1011011011 : tanh_out_reg <= 10'b1100110000;
		12'b1011011100 : tanh_out_reg <= 10'b1100110000;
		12'b1011011101 : tanh_out_reg <= 10'b1100110000;
		12'b1011011110 : tanh_out_reg <= 10'b1100110001;
		12'b1011011111 : tanh_out_reg <= 10'b1100110001;
		12'b1011100000 : tanh_out_reg <= 10'b1100110001;
		12'b1011100001 : tanh_out_reg <= 10'b1100110010;
		12'b1011100010 : tanh_out_reg <= 10'b1100110010;
		12'b1011100011 : tanh_out_reg <= 10'b1100110010;
		12'b1011100100 : tanh_out_reg <= 10'b1100110011;
		12'b1011100101 : tanh_out_reg <= 10'b1100110011;
		12'b1011100110 : tanh_out_reg <= 10'b1100110011;
		12'b1011100111 : tanh_out_reg <= 10'b1100110100;
		12'b1011101000 : tanh_out_reg <= 10'b1100110100;
		12'b1011101001 : tanh_out_reg <= 10'b1100110101;
		12'b1011101010 : tanh_out_reg <= 10'b1100110101;
		12'b1011101011 : tanh_out_reg <= 10'b1100110101;
		12'b1011101100 : tanh_out_reg <= 10'b1100110110;
		12'b1011101101 : tanh_out_reg <= 10'b1100110110;
		12'b1011101110 : tanh_out_reg <= 10'b1100110110;
		12'b1011101111 : tanh_out_reg <= 10'b1100110111;
		12'b1011110000 : tanh_out_reg <= 10'b1100110111;
		12'b1011110001 : tanh_out_reg <= 10'b1100111000;
		12'b1011110010 : tanh_out_reg <= 10'b1100111000;
		12'b1011110011 : tanh_out_reg <= 10'b1100111000;
		12'b1011110100 : tanh_out_reg <= 10'b1100111001;
		12'b1011110101 : tanh_out_reg <= 10'b1100111001;
		12'b1011110110 : tanh_out_reg <= 10'b1100111001;
		12'b1011110111 : tanh_out_reg <= 10'b1100111010;
		12'b1011111000 : tanh_out_reg <= 10'b1100111010;
		12'b1011111001 : tanh_out_reg <= 10'b1100111011;
		12'b1011111010 : tanh_out_reg <= 10'b1100111011;
		12'b1011111011 : tanh_out_reg <= 10'b1100111011;
		12'b1011111100 : tanh_out_reg <= 10'b1100111100;
		12'b1011111101 : tanh_out_reg <= 10'b1100111100;
		12'b1011111110 : tanh_out_reg <= 10'b1100111101;
		12'b1011111111 : tanh_out_reg <= 10'b1100111101;
		12'b1100000000 : tanh_out_reg <= 10'b1100111110;
		12'b1100000001 : tanh_out_reg <= 10'b1100111110;
		12'b1100000010 : tanh_out_reg <= 10'b1100111110;
		12'b1100000011 : tanh_out_reg <= 10'b1100111111;
		12'b1100000100 : tanh_out_reg <= 10'b1100111111;
		12'b1100000101 : tanh_out_reg <= 10'b1101000000;
		12'b1100000110 : tanh_out_reg <= 10'b1101000000;
		12'b1100000111 : tanh_out_reg <= 10'b1101000001;
		12'b1100001000 : tanh_out_reg <= 10'b1101000001;
		12'b1100001001 : tanh_out_reg <= 10'b1101000001;
		12'b1100001010 : tanh_out_reg <= 10'b1101000010;
		12'b1100001011 : tanh_out_reg <= 10'b1101000010;
		12'b1100001100 : tanh_out_reg <= 10'b1101000011;
		12'b1100001101 : tanh_out_reg <= 10'b1101000011;
		12'b1100001110 : tanh_out_reg <= 10'b1101000100;
		12'b1100001111 : tanh_out_reg <= 10'b1101000100;
		12'b1100010000 : tanh_out_reg <= 10'b1101000101;
		12'b1100010001 : tanh_out_reg <= 10'b1101000101;
		12'b1100010010 : tanh_out_reg <= 10'b1101000110;
		12'b1100010011 : tanh_out_reg <= 10'b1101000110;
		12'b1100010100 : tanh_out_reg <= 10'b1101000110;
		12'b1100010101 : tanh_out_reg <= 10'b1101000111;
		12'b1100010110 : tanh_out_reg <= 10'b1101000111;
		12'b1100010111 : tanh_out_reg <= 10'b1101001000;
		12'b1100011000 : tanh_out_reg <= 10'b1101001000;
		12'b1100011001 : tanh_out_reg <= 10'b1101001001;
		12'b1100011010 : tanh_out_reg <= 10'b1101001001;
		12'b1100011011 : tanh_out_reg <= 10'b1101001010;
		12'b1100011100 : tanh_out_reg <= 10'b1101001010;
		12'b1100011101 : tanh_out_reg <= 10'b1101001011;
		12'b1100011110 : tanh_out_reg <= 10'b1101001011;
		12'b1100011111 : tanh_out_reg <= 10'b1101001100;
		12'b1100100000 : tanh_out_reg <= 10'b1101001100;
		12'b1100100001 : tanh_out_reg <= 10'b1101001101;
		12'b1100100010 : tanh_out_reg <= 10'b1101001101;
		12'b1100100011 : tanh_out_reg <= 10'b1101001110;
		12'b1100100100 : tanh_out_reg <= 10'b1101001110;
		12'b1100100101 : tanh_out_reg <= 10'b1101001111;
		12'b1100100110 : tanh_out_reg <= 10'b1101001111;
		12'b1100100111 : tanh_out_reg <= 10'b1101010000;
		12'b1100101000 : tanh_out_reg <= 10'b1101010000;
		12'b1100101001 : tanh_out_reg <= 10'b1101010001;
		12'b1100101010 : tanh_out_reg <= 10'b1101010001;
		12'b1100101011 : tanh_out_reg <= 10'b1101010010;
		12'b1100101100 : tanh_out_reg <= 10'b1101010011;
		12'b1100101101 : tanh_out_reg <= 10'b1101010011;
		12'b1100101110 : tanh_out_reg <= 10'b1101010100;
		12'b1100101111 : tanh_out_reg <= 10'b1101010100;
		12'b1100110000 : tanh_out_reg <= 10'b1101010101;
		12'b1100110001 : tanh_out_reg <= 10'b1101010101;
		12'b1100110010 : tanh_out_reg <= 10'b1101010110;
		12'b1100110011 : tanh_out_reg <= 10'b1101010110;
		12'b1100110100 : tanh_out_reg <= 10'b1101010111;
		12'b1100110101 : tanh_out_reg <= 10'b1101011000;
		12'b1100110110 : tanh_out_reg <= 10'b1101011000;
		12'b1100110111 : tanh_out_reg <= 10'b1101011001;
		12'b1100111000 : tanh_out_reg <= 10'b1101011001;
		12'b1100111001 : tanh_out_reg <= 10'b1101011010;
		12'b1100111010 : tanh_out_reg <= 10'b1101011010;
		12'b1100111011 : tanh_out_reg <= 10'b1101011011;
		12'b1100111100 : tanh_out_reg <= 10'b1101011100;
		12'b1100111101 : tanh_out_reg <= 10'b1101011100;
		12'b1100111110 : tanh_out_reg <= 10'b1101011101;
		12'b1100111111 : tanh_out_reg <= 10'b1101011101;
		12'b1101000000 : tanh_out_reg <= 10'b1101011110;
		12'b1101000001 : tanh_out_reg <= 10'b1101011110;
		12'b1101000010 : tanh_out_reg <= 10'b1101011111;
		12'b1101000011 : tanh_out_reg <= 10'b1101100000;
		12'b1101000100 : tanh_out_reg <= 10'b1101100000;
		12'b1101000101 : tanh_out_reg <= 10'b1101100001;
		12'b1101000110 : tanh_out_reg <= 10'b1101100010;
		12'b1101000111 : tanh_out_reg <= 10'b1101100010;
		12'b1101001000 : tanh_out_reg <= 10'b1101100011;
		12'b1101001001 : tanh_out_reg <= 10'b1101100011;
		12'b1101001010 : tanh_out_reg <= 10'b1101100100;
		12'b1101001011 : tanh_out_reg <= 10'b1101100101;
		12'b1101001100 : tanh_out_reg <= 10'b1101100101;
		12'b1101001101 : tanh_out_reg <= 10'b1101100110;
		12'b1101001110 : tanh_out_reg <= 10'b1101100111;
		12'b1101001111 : tanh_out_reg <= 10'b1101100111;
		12'b1101010000 : tanh_out_reg <= 10'b1101101000;
		12'b1101010001 : tanh_out_reg <= 10'b1101101000;
		12'b1101010010 : tanh_out_reg <= 10'b1101101001;
		12'b1101010011 : tanh_out_reg <= 10'b1101101010;
		12'b1101010100 : tanh_out_reg <= 10'b1101101010;
		12'b1101010101 : tanh_out_reg <= 10'b1101101011;
		12'b1101010110 : tanh_out_reg <= 10'b1101101100;
		12'b1101010111 : tanh_out_reg <= 10'b1101101100;
		12'b1101011000 : tanh_out_reg <= 10'b1101101101;
		12'b1101011001 : tanh_out_reg <= 10'b1101101110;
		12'b1101011010 : tanh_out_reg <= 10'b1101101110;
		12'b1101011011 : tanh_out_reg <= 10'b1101101111;
		12'b1101011100 : tanh_out_reg <= 10'b1101110000;
		12'b1101011101 : tanh_out_reg <= 10'b1101110000;
		12'b1101011110 : tanh_out_reg <= 10'b1101110001;
		12'b1101011111 : tanh_out_reg <= 10'b1101110010;
		12'b1101100000 : tanh_out_reg <= 10'b1101110011;
		12'b1101100001 : tanh_out_reg <= 10'b1101110011;
		12'b1101100010 : tanh_out_reg <= 10'b1101110100;
		12'b1101100011 : tanh_out_reg <= 10'b1101110101;
		12'b1101100100 : tanh_out_reg <= 10'b1101110101;
		12'b1101100101 : tanh_out_reg <= 10'b1101110110;
		12'b1101100110 : tanh_out_reg <= 10'b1101110111;
		12'b1101100111 : tanh_out_reg <= 10'b1101110111;
		12'b1101101000 : tanh_out_reg <= 10'b1101111000;
		12'b1101101001 : tanh_out_reg <= 10'b1101111001;
		12'b1101101010 : tanh_out_reg <= 10'b1101111010;
		12'b1101101011 : tanh_out_reg <= 10'b1101111010;
		12'b1101101100 : tanh_out_reg <= 10'b1101111011;
		12'b1101101101 : tanh_out_reg <= 10'b1101111100;
		12'b1101101110 : tanh_out_reg <= 10'b1101111101;
		12'b1101101111 : tanh_out_reg <= 10'b1101111101;
		12'b1101110000 : tanh_out_reg <= 10'b1101111110;
		12'b1101110001 : tanh_out_reg <= 10'b1101111111;
		12'b1101110010 : tanh_out_reg <= 10'b1101111111;
		12'b1101110011 : tanh_out_reg <= 10'b1110000000;
		12'b1101110100 : tanh_out_reg <= 10'b1110000001;
		12'b1101110101 : tanh_out_reg <= 10'b1110000010;
		12'b1101110110 : tanh_out_reg <= 10'b1110000010;
		12'b1101110111 : tanh_out_reg <= 10'b1110000011;
		12'b1101111000 : tanh_out_reg <= 10'b1110000100;
		12'b1101111001 : tanh_out_reg <= 10'b1110000101;
		12'b1101111010 : tanh_out_reg <= 10'b1110000110;
		12'b1101111011 : tanh_out_reg <= 10'b1110000110;
		12'b1101111100 : tanh_out_reg <= 10'b1110000111;
		12'b1101111101 : tanh_out_reg <= 10'b1110001000;
		12'b1101111110 : tanh_out_reg <= 10'b1110001001;
		12'b1101111111 : tanh_out_reg <= 10'b1110001001;
		12'b1110000000 : tanh_out_reg <= 10'b1110001010;
		12'b1110000001 : tanh_out_reg <= 10'b1110001011;
		12'b1110000010 : tanh_out_reg <= 10'b1110001100;
		12'b1110000011 : tanh_out_reg <= 10'b1110001101;
		12'b1110000100 : tanh_out_reg <= 10'b1110001101;
		12'b1110000101 : tanh_out_reg <= 10'b1110001110;
		12'b1110000110 : tanh_out_reg <= 10'b1110001111;
		12'b1110000111 : tanh_out_reg <= 10'b1110010000;
		12'b1110001000 : tanh_out_reg <= 10'b1110010001;
		12'b1110001001 : tanh_out_reg <= 10'b1110010001;
		12'b1110001010 : tanh_out_reg <= 10'b1110010010;
		12'b1110001011 : tanh_out_reg <= 10'b1110010011;
		12'b1110001100 : tanh_out_reg <= 10'b1110010100;
		12'b1110001101 : tanh_out_reg <= 10'b1110010101;
		12'b1110001110 : tanh_out_reg <= 10'b1110010101;
		12'b1110001111 : tanh_out_reg <= 10'b1110010110;
		12'b1110010000 : tanh_out_reg <= 10'b1110010111;
		12'b1110010001 : tanh_out_reg <= 10'b1110011000;
		12'b1110010010 : tanh_out_reg <= 10'b1110011001;
		12'b1110010011 : tanh_out_reg <= 10'b1110011010;
		12'b1110010100 : tanh_out_reg <= 10'b1110011010;
		12'b1110010101 : tanh_out_reg <= 10'b1110011011;
		12'b1110010110 : tanh_out_reg <= 10'b1110011100;
		12'b1110010111 : tanh_out_reg <= 10'b1110011101;
		12'b1110011000 : tanh_out_reg <= 10'b1110011110;
		12'b1110011001 : tanh_out_reg <= 10'b1110011111;
		12'b1110011010 : tanh_out_reg <= 10'b1110100000;
		12'b1110011011 : tanh_out_reg <= 10'b1110100000;
		12'b1110011100 : tanh_out_reg <= 10'b1110100001;
		12'b1110011101 : tanh_out_reg <= 10'b1110100010;
		12'b1110011110 : tanh_out_reg <= 10'b1110100011;
		12'b1110011111 : tanh_out_reg <= 10'b1110100100;
		12'b1110100000 : tanh_out_reg <= 10'b1110100101;
		12'b1110100001 : tanh_out_reg <= 10'b1110100110;
		12'b1110100010 : tanh_out_reg <= 10'b1110100111;
		12'b1110100011 : tanh_out_reg <= 10'b1110100111;
		12'b1110100100 : tanh_out_reg <= 10'b1110101000;
		12'b1110100101 : tanh_out_reg <= 10'b1110101001;
		12'b1110100110 : tanh_out_reg <= 10'b1110101010;
		12'b1110100111 : tanh_out_reg <= 10'b1110101011;
		12'b1110101000 : tanh_out_reg <= 10'b1110101100;
		12'b1110101001 : tanh_out_reg <= 10'b1110101101;
		12'b1110101010 : tanh_out_reg <= 10'b1110101110;
		12'b1110101011 : tanh_out_reg <= 10'b1110101110;
		12'b1110101100 : tanh_out_reg <= 10'b1110101111;
		12'b1110101101 : tanh_out_reg <= 10'b1110110000;
		12'b1110101110 : tanh_out_reg <= 10'b1110110001;
		12'b1110101111 : tanh_out_reg <= 10'b1110110010;
		12'b1110110000 : tanh_out_reg <= 10'b1110110011;
		12'b1110110001 : tanh_out_reg <= 10'b1110110100;
		12'b1110110010 : tanh_out_reg <= 10'b1110110101;
		12'b1110110011 : tanh_out_reg <= 10'b1110110110;
		12'b1110110100 : tanh_out_reg <= 10'b1110110111;
		12'b1110110101 : tanh_out_reg <= 10'b1110111000;
		12'b1110110110 : tanh_out_reg <= 10'b1110111000;
		12'b1110110111 : tanh_out_reg <= 10'b1110111001;
		12'b1110111000 : tanh_out_reg <= 10'b1110111010;
		12'b1110111001 : tanh_out_reg <= 10'b1110111011;
		12'b1110111010 : tanh_out_reg <= 10'b1110111100;
		12'b1110111011 : tanh_out_reg <= 10'b1110111101;
		12'b1110111100 : tanh_out_reg <= 10'b1110111110;
		12'b1110111101 : tanh_out_reg <= 10'b1110111111;
		12'b1110111110 : tanh_out_reg <= 10'b1111000000;
		12'b1110111111 : tanh_out_reg <= 10'b1111000001;
		12'b1111000000 : tanh_out_reg <= 10'b1111000010;
		12'b1111000001 : tanh_out_reg <= 10'b1111000011;
		12'b1111000010 : tanh_out_reg <= 10'b1111000100;
		12'b1111000011 : tanh_out_reg <= 10'b1111000101;
		12'b1111000100 : tanh_out_reg <= 10'b1111000110;
		12'b1111000101 : tanh_out_reg <= 10'b1111000111;
		12'b1111000110 : tanh_out_reg <= 10'b1111000111;
		12'b1111000111 : tanh_out_reg <= 10'b1111001000;
		12'b1111001000 : tanh_out_reg <= 10'b1111001001;
		12'b1111001001 : tanh_out_reg <= 10'b1111001010;
		12'b1111001010 : tanh_out_reg <= 10'b1111001011;
		12'b1111001011 : tanh_out_reg <= 10'b1111001100;
		12'b1111001100 : tanh_out_reg <= 10'b1111001101;
		12'b1111001101 : tanh_out_reg <= 10'b1111001110;
		12'b1111001110 : tanh_out_reg <= 10'b1111001111;
		12'b1111001111 : tanh_out_reg <= 10'b1111010000;
		12'b1111010000 : tanh_out_reg <= 10'b1111010001;
		12'b1111010001 : tanh_out_reg <= 10'b1111010010;
		12'b1111010010 : tanh_out_reg <= 10'b1111010011;
		12'b1111010011 : tanh_out_reg <= 10'b1111010100;
		12'b1111010100 : tanh_out_reg <= 10'b1111010101;
		12'b1111010101 : tanh_out_reg <= 10'b1111010110;
		12'b1111010110 : tanh_out_reg <= 10'b1111010111;
		12'b1111010111 : tanh_out_reg <= 10'b1111011000;
		12'b1111011000 : tanh_out_reg <= 10'b1111011001;
		12'b1111011001 : tanh_out_reg <= 10'b1111011010;
		12'b1111011010 : tanh_out_reg <= 10'b1111011011;
		12'b1111011011 : tanh_out_reg <= 10'b1111011100;
		12'b1111011100 : tanh_out_reg <= 10'b1111011101;
		12'b1111011101 : tanh_out_reg <= 10'b1111011110;
		12'b1111011110 : tanh_out_reg <= 10'b1111011111;
		12'b1111011111 : tanh_out_reg <= 10'b1111100000;
		12'b1111100000 : tanh_out_reg <= 10'b1111100001;
		12'b1111100001 : tanh_out_reg <= 10'b1111100010;
		12'b1111100010 : tanh_out_reg <= 10'b1111100011;
		12'b1111100011 : tanh_out_reg <= 10'b1111100100;
		12'b1111100100 : tanh_out_reg <= 10'b1111100101;
		12'b1111100101 : tanh_out_reg <= 10'b1111100110;
		12'b1111100110 : tanh_out_reg <= 10'b1111100111;
		12'b1111100111 : tanh_out_reg <= 10'b1111101000;
		12'b1111101000 : tanh_out_reg <= 10'b1111101001;
		12'b1111101001 : tanh_out_reg <= 10'b1111101010;
		12'b1111101010 : tanh_out_reg <= 10'b1111101011;
		12'b1111101011 : tanh_out_reg <= 10'b1111101100;
		12'b1111101100 : tanh_out_reg <= 10'b1111101101;
		12'b1111101101 : tanh_out_reg <= 10'b1111101110;
		12'b1111101110 : tanh_out_reg <= 10'b1111101111;
		12'b1111101111 : tanh_out_reg <= 10'b1111110000;
		12'b1111110000 : tanh_out_reg <= 10'b1111110001;
		12'b1111110001 : tanh_out_reg <= 10'b1111110010;
		12'b1111110010 : tanh_out_reg <= 10'b1111110011;
		12'b1111110011 : tanh_out_reg <= 10'b1111110100;
		12'b1111110100 : tanh_out_reg <= 10'b1111110101;
		12'b1111110101 : tanh_out_reg <= 10'b1111110110;
		12'b1111110110 : tanh_out_reg <= 10'b1111110111;
		12'b1111110111 : tanh_out_reg <= 10'b1111111000;
		12'b1111111000 : tanh_out_reg <= 10'b1111111001;
		12'b1111111001 : tanh_out_reg <= 10'b1111111010;
		12'b1111111010 : tanh_out_reg <= 10'b1111111011;
		12'b1111111011 : tanh_out_reg <= 10'b1111111100;
		12'b1111111100 : tanh_out_reg <= 10'b1111111101;
		12'b1111111101 : tanh_out_reg <= 10'b1111111110;
		12'b1111111110 : tanh_out_reg <= 10'b1111111111;
		12'b1111111111 : tanh_out_reg <= 10'b0000000000;
	endcase
end

endmodule
