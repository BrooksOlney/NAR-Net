`timescale 1ns / 1ps
module tanh_lut #(parameter N=8, parameter Q=7) (
	input [N-1:0] addr,
	 input clk,
	 output signed [N-1:0] tanh_out
	);
reg signed [N-1:0] tanh_out_reg;
assign tanh_out = tanh_out_reg;

always @(negedge clk) begin
	case (addr)
		12'b00000000 : tanh_out_reg <= 8'b00000000;
		12'b00000001 : tanh_out_reg <= 8'b00000000;
		12'b00000010 : tanh_out_reg <= 8'b00000001;
		12'b00000011 : tanh_out_reg <= 8'b00000010;
		12'b00000100 : tanh_out_reg <= 8'b00000011;
		12'b00000101 : tanh_out_reg <= 8'b00000100;
		12'b00000110 : tanh_out_reg <= 8'b00000101;
		12'b00000111 : tanh_out_reg <= 8'b00000110;
		12'b00001000 : tanh_out_reg <= 8'b00000111;
		12'b00001001 : tanh_out_reg <= 8'b00001000;
		12'b00001010 : tanh_out_reg <= 8'b00001001;
		12'b00001011 : tanh_out_reg <= 8'b00001010;
		12'b00001100 : tanh_out_reg <= 8'b00001011;
		12'b00001101 : tanh_out_reg <= 8'b00001100;
		12'b00001110 : tanh_out_reg <= 8'b00001101;
		12'b00001111 : tanh_out_reg <= 8'b00001110;
		12'b00010000 : tanh_out_reg <= 8'b00001111;
		12'b00010001 : tanh_out_reg <= 8'b00010000;
		12'b00010010 : tanh_out_reg <= 8'b00010001;
		12'b00010011 : tanh_out_reg <= 8'b00010010;
		12'b00010100 : tanh_out_reg <= 8'b00010011;
		12'b00010101 : tanh_out_reg <= 8'b00010100;
		12'b00010110 : tanh_out_reg <= 8'b00010101;
		12'b00010111 : tanh_out_reg <= 8'b00010110;
		12'b00011000 : tanh_out_reg <= 8'b00010111;
		12'b00011001 : tanh_out_reg <= 8'b00011000;
		12'b00011010 : tanh_out_reg <= 8'b00011001;
		12'b00011011 : tanh_out_reg <= 8'b00011010;
		12'b00011100 : tanh_out_reg <= 8'b00011011;
		12'b00011101 : tanh_out_reg <= 8'b00011100;
		12'b00011110 : tanh_out_reg <= 8'b00011101;
		12'b00011111 : tanh_out_reg <= 8'b00011110;
		12'b00100000 : tanh_out_reg <= 8'b00011111;
		12'b00100001 : tanh_out_reg <= 8'b00100000;
		12'b00100010 : tanh_out_reg <= 8'b00100001;
		12'b00100011 : tanh_out_reg <= 8'b00100010;
		12'b00100100 : tanh_out_reg <= 8'b00100011;
		12'b00100101 : tanh_out_reg <= 8'b00100100;
		12'b00100110 : tanh_out_reg <= 8'b00100100;
		12'b00100111 : tanh_out_reg <= 8'b00100101;
		12'b00101000 : tanh_out_reg <= 8'b00100110;
		12'b00101001 : tanh_out_reg <= 8'b00100111;
		12'b00101010 : tanh_out_reg <= 8'b00101000;
		12'b00101011 : tanh_out_reg <= 8'b00101001;
		12'b00101100 : tanh_out_reg <= 8'b00101010;
		12'b00101101 : tanh_out_reg <= 8'b00101011;
		12'b00101110 : tanh_out_reg <= 8'b00101100;
		12'b00101111 : tanh_out_reg <= 8'b00101100;
		12'b00110000 : tanh_out_reg <= 8'b00101101;
		12'b00110001 : tanh_out_reg <= 8'b00101110;
		12'b00110010 : tanh_out_reg <= 8'b00101111;
		12'b00110011 : tanh_out_reg <= 8'b00110000;
		12'b00110100 : tanh_out_reg <= 8'b00110001;
		12'b00110101 : tanh_out_reg <= 8'b00110010;
		12'b00110110 : tanh_out_reg <= 8'b00110011;
		12'b00110111 : tanh_out_reg <= 8'b00110011;
		12'b00111000 : tanh_out_reg <= 8'b00110100;
		12'b00111001 : tanh_out_reg <= 8'b00110101;
		12'b00111010 : tanh_out_reg <= 8'b00110110;
		12'b00111011 : tanh_out_reg <= 8'b00110111;
		12'b00111100 : tanh_out_reg <= 8'b00110111;
		12'b00111101 : tanh_out_reg <= 8'b00111000;
		12'b00111110 : tanh_out_reg <= 8'b00111001;
		12'b00111111 : tanh_out_reg <= 8'b00111010;
		12'b01000000 : tanh_out_reg <= 8'b00111011;
		12'b01000001 : tanh_out_reg <= 8'b00111011;
		12'b01000010 : tanh_out_reg <= 8'b00111100;
		12'b01000011 : tanh_out_reg <= 8'b00111101;
		12'b01000100 : tanh_out_reg <= 8'b00111110;
		12'b01000101 : tanh_out_reg <= 8'b00111111;
		12'b01000110 : tanh_out_reg <= 8'b00111111;
		12'b01000111 : tanh_out_reg <= 8'b01000000;
		12'b01001000 : tanh_out_reg <= 8'b01000001;
		12'b01001001 : tanh_out_reg <= 8'b01000001;
		12'b01001010 : tanh_out_reg <= 8'b01000010;
		12'b01001011 : tanh_out_reg <= 8'b01000011;
		12'b01001100 : tanh_out_reg <= 8'b01000100;
		12'b01001101 : tanh_out_reg <= 8'b01000100;
		12'b01001110 : tanh_out_reg <= 8'b01000101;
		12'b01001111 : tanh_out_reg <= 8'b01000110;
		12'b01010000 : tanh_out_reg <= 8'b01000110;
		12'b01010001 : tanh_out_reg <= 8'b01000111;
		12'b01010010 : tanh_out_reg <= 8'b01001000;
		12'b01010011 : tanh_out_reg <= 8'b01001001;
		12'b01010100 : tanh_out_reg <= 8'b01001001;
		12'b01010101 : tanh_out_reg <= 8'b01001010;
		12'b01010110 : tanh_out_reg <= 8'b01001011;
		12'b01010111 : tanh_out_reg <= 8'b01001011;
		12'b01011000 : tanh_out_reg <= 8'b01001100;
		12'b01011001 : tanh_out_reg <= 8'b01001100;
		12'b01011010 : tanh_out_reg <= 8'b01001101;
		12'b01011011 : tanh_out_reg <= 8'b01001110;
		12'b01011100 : tanh_out_reg <= 8'b01001110;
		12'b01011101 : tanh_out_reg <= 8'b01001111;
		12'b01011110 : tanh_out_reg <= 8'b01010000;
		12'b01011111 : tanh_out_reg <= 8'b01010000;
		12'b01100000 : tanh_out_reg <= 8'b01010001;
		12'b01100001 : tanh_out_reg <= 8'b01010001;
		12'b01100010 : tanh_out_reg <= 8'b01010010;
		12'b01100011 : tanh_out_reg <= 8'b01010011;
		12'b01100100 : tanh_out_reg <= 8'b01010011;
		12'b01100101 : tanh_out_reg <= 8'b01010100;
		12'b01100110 : tanh_out_reg <= 8'b01010100;
		12'b01100111 : tanh_out_reg <= 8'b01010101;
		12'b01101000 : tanh_out_reg <= 8'b01010101;
		12'b01101001 : tanh_out_reg <= 8'b01010110;
		12'b01101010 : tanh_out_reg <= 8'b01010110;
		12'b01101011 : tanh_out_reg <= 8'b01010111;
		12'b01101100 : tanh_out_reg <= 8'b01011000;
		12'b01101101 : tanh_out_reg <= 8'b01011000;
		12'b01101110 : tanh_out_reg <= 8'b01011001;
		12'b01101111 : tanh_out_reg <= 8'b01011001;
		12'b01110000 : tanh_out_reg <= 8'b01011010;
		12'b01110001 : tanh_out_reg <= 8'b01011010;
		12'b01110010 : tanh_out_reg <= 8'b01011011;
		12'b01110011 : tanh_out_reg <= 8'b01011011;
		12'b01110100 : tanh_out_reg <= 8'b01011100;
		12'b01110101 : tanh_out_reg <= 8'b01011100;
		12'b01110110 : tanh_out_reg <= 8'b01011101;
		12'b01110111 : tanh_out_reg <= 8'b01011101;
		12'b01111000 : tanh_out_reg <= 8'b01011101;
		12'b01111001 : tanh_out_reg <= 8'b01011110;
		12'b01111010 : tanh_out_reg <= 8'b01011110;
		12'b01111011 : tanh_out_reg <= 8'b01011111;
		12'b01111100 : tanh_out_reg <= 8'b01011111;
		12'b01111101 : tanh_out_reg <= 8'b01100000;
		12'b01111110 : tanh_out_reg <= 8'b01100000;
		12'b01111111 : tanh_out_reg <= 8'b01100001;
		12'b10000000 : tanh_out_reg <= 8'b10011111;
		12'b10000001 : tanh_out_reg <= 8'b10011111;
		12'b10000010 : tanh_out_reg <= 8'b10100000;
		12'b10000011 : tanh_out_reg <= 8'b10100000;
		12'b10000100 : tanh_out_reg <= 8'b10100001;
		12'b10000101 : tanh_out_reg <= 8'b10100001;
		12'b10000110 : tanh_out_reg <= 8'b10100010;
		12'b10000111 : tanh_out_reg <= 8'b10100010;
		12'b10001000 : tanh_out_reg <= 8'b10100011;
		12'b10001001 : tanh_out_reg <= 8'b10100011;
		12'b10001010 : tanh_out_reg <= 8'b10100011;
		12'b10001011 : tanh_out_reg <= 8'b10100100;
		12'b10001100 : tanh_out_reg <= 8'b10100100;
		12'b10001101 : tanh_out_reg <= 8'b10100101;
		12'b10001110 : tanh_out_reg <= 8'b10100101;
		12'b10001111 : tanh_out_reg <= 8'b10100110;
		12'b10010000 : tanh_out_reg <= 8'b10100110;
		12'b10010001 : tanh_out_reg <= 8'b10100111;
		12'b10010010 : tanh_out_reg <= 8'b10100111;
		12'b10010011 : tanh_out_reg <= 8'b10101000;
		12'b10010100 : tanh_out_reg <= 8'b10101000;
		12'b10010101 : tanh_out_reg <= 8'b10101001;
		12'b10010110 : tanh_out_reg <= 8'b10101010;
		12'b10010111 : tanh_out_reg <= 8'b10101010;
		12'b10011000 : tanh_out_reg <= 8'b10101011;
		12'b10011001 : tanh_out_reg <= 8'b10101011;
		12'b10011010 : tanh_out_reg <= 8'b10101100;
		12'b10011011 : tanh_out_reg <= 8'b10101100;
		12'b10011100 : tanh_out_reg <= 8'b10101101;
		12'b10011101 : tanh_out_reg <= 8'b10101101;
		12'b10011110 : tanh_out_reg <= 8'b10101110;
		12'b10011111 : tanh_out_reg <= 8'b10101111;
		12'b10100000 : tanh_out_reg <= 8'b10101111;
		12'b10100001 : tanh_out_reg <= 8'b10110000;
		12'b10100010 : tanh_out_reg <= 8'b10110000;
		12'b10100011 : tanh_out_reg <= 8'b10110001;
		12'b10100100 : tanh_out_reg <= 8'b10110010;
		12'b10100101 : tanh_out_reg <= 8'b10110010;
		12'b10100110 : tanh_out_reg <= 8'b10110011;
		12'b10100111 : tanh_out_reg <= 8'b10110100;
		12'b10101000 : tanh_out_reg <= 8'b10110100;
		12'b10101001 : tanh_out_reg <= 8'b10110101;
		12'b10101010 : tanh_out_reg <= 8'b10110101;
		12'b10101011 : tanh_out_reg <= 8'b10110110;
		12'b10101100 : tanh_out_reg <= 8'b10110111;
		12'b10101101 : tanh_out_reg <= 8'b10110111;
		12'b10101110 : tanh_out_reg <= 8'b10111000;
		12'b10101111 : tanh_out_reg <= 8'b10111001;
		12'b10110000 : tanh_out_reg <= 8'b10111010;
		12'b10110001 : tanh_out_reg <= 8'b10111010;
		12'b10110010 : tanh_out_reg <= 8'b10111011;
		12'b10110011 : tanh_out_reg <= 8'b10111100;
		12'b10110100 : tanh_out_reg <= 8'b10111100;
		12'b10110101 : tanh_out_reg <= 8'b10111101;
		12'b10110110 : tanh_out_reg <= 8'b10111110;
		12'b10110111 : tanh_out_reg <= 8'b10111111;
		12'b10111000 : tanh_out_reg <= 8'b10111111;
		12'b10111001 : tanh_out_reg <= 8'b11000000;
		12'b10111010 : tanh_out_reg <= 8'b11000001;
		12'b10111011 : tanh_out_reg <= 8'b11000001;
		12'b10111100 : tanh_out_reg <= 8'b11000010;
		12'b10111101 : tanh_out_reg <= 8'b11000011;
		12'b10111110 : tanh_out_reg <= 8'b11000100;
		12'b10111111 : tanh_out_reg <= 8'b11000101;
		12'b11000000 : tanh_out_reg <= 8'b11000101;
		12'b11000001 : tanh_out_reg <= 8'b11000110;
		12'b11000010 : tanh_out_reg <= 8'b11000111;
		12'b11000011 : tanh_out_reg <= 8'b11001000;
		12'b11000100 : tanh_out_reg <= 8'b11001001;
		12'b11000101 : tanh_out_reg <= 8'b11001001;
		12'b11000110 : tanh_out_reg <= 8'b11001010;
		12'b11000111 : tanh_out_reg <= 8'b11001011;
		12'b11001000 : tanh_out_reg <= 8'b11001100;
		12'b11001001 : tanh_out_reg <= 8'b11001101;
		12'b11001010 : tanh_out_reg <= 8'b11001101;
		12'b11001011 : tanh_out_reg <= 8'b11001110;
		12'b11001100 : tanh_out_reg <= 8'b11001111;
		12'b11001101 : tanh_out_reg <= 8'b11010000;
		12'b11001110 : tanh_out_reg <= 8'b11010001;
		12'b11001111 : tanh_out_reg <= 8'b11010010;
		12'b11010000 : tanh_out_reg <= 8'b11010011;
		12'b11010001 : tanh_out_reg <= 8'b11010100;
		12'b11010010 : tanh_out_reg <= 8'b11010100;
		12'b11010011 : tanh_out_reg <= 8'b11010101;
		12'b11010100 : tanh_out_reg <= 8'b11010110;
		12'b11010101 : tanh_out_reg <= 8'b11010111;
		12'b11010110 : tanh_out_reg <= 8'b11011000;
		12'b11010111 : tanh_out_reg <= 8'b11011001;
		12'b11011000 : tanh_out_reg <= 8'b11011010;
		12'b11011001 : tanh_out_reg <= 8'b11011011;
		12'b11011010 : tanh_out_reg <= 8'b11011100;
		12'b11011011 : tanh_out_reg <= 8'b11011100;
		12'b11011100 : tanh_out_reg <= 8'b11011101;
		12'b11011101 : tanh_out_reg <= 8'b11011110;
		12'b11011110 : tanh_out_reg <= 8'b11011111;
		12'b11011111 : tanh_out_reg <= 8'b11100000;
		12'b11100000 : tanh_out_reg <= 8'b11100001;
		12'b11100001 : tanh_out_reg <= 8'b11100010;
		12'b11100010 : tanh_out_reg <= 8'b11100011;
		12'b11100011 : tanh_out_reg <= 8'b11100100;
		12'b11100100 : tanh_out_reg <= 8'b11100101;
		12'b11100101 : tanh_out_reg <= 8'b11100110;
		12'b11100110 : tanh_out_reg <= 8'b11100111;
		12'b11100111 : tanh_out_reg <= 8'b11101000;
		12'b11101000 : tanh_out_reg <= 8'b11101001;
		12'b11101001 : tanh_out_reg <= 8'b11101010;
		12'b11101010 : tanh_out_reg <= 8'b11101011;
		12'b11101011 : tanh_out_reg <= 8'b11101100;
		12'b11101100 : tanh_out_reg <= 8'b11101101;
		12'b11101101 : tanh_out_reg <= 8'b11101110;
		12'b11101110 : tanh_out_reg <= 8'b11101111;
		12'b11101111 : tanh_out_reg <= 8'b11110000;
		12'b11110000 : tanh_out_reg <= 8'b11110001;
		12'b11110001 : tanh_out_reg <= 8'b11110010;
		12'b11110010 : tanh_out_reg <= 8'b11110011;
		12'b11110011 : tanh_out_reg <= 8'b11110100;
		12'b11110100 : tanh_out_reg <= 8'b11110101;
		12'b11110101 : tanh_out_reg <= 8'b11110110;
		12'b11110110 : tanh_out_reg <= 8'b11110111;
		12'b11110111 : tanh_out_reg <= 8'b11111000;
		12'b11111000 : tanh_out_reg <= 8'b11111001;
		12'b11111001 : tanh_out_reg <= 8'b11111010;
		12'b11111010 : tanh_out_reg <= 8'b11111011;
		12'b11111011 : tanh_out_reg <= 8'b11111100;
		12'b11111100 : tanh_out_reg <= 8'b11111101;
		12'b11111101 : tanh_out_reg <= 8'b11111110;
		12'b11111110 : tanh_out_reg <= 8'b11111111;
		12'b11111111 : tanh_out_reg <= 8'b00000000;
	endcase
end

endmodule
